module (input clk, input rst, input N, output reg F);

    
    always @ (posedge clk) begin
        if 
    end
    

endmodule
